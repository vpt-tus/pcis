package bcd;
	typedef logic [3:0] bcd_t;
endpackage