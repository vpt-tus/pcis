import bcd::*;

module bcd_adder_1d(
  input bcd_t a,b,
  input cin,
  output bcd_t s,
  output logic cout);

  // TODO
  
endmodule