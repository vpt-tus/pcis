import bcd::*;

module bcd_adder_3d(
	input bcd_t [2:0] op1, op2,
	input cin,
	output bcd_t [2:0] sum,
	output logic cout);

	// TODO

endmodule