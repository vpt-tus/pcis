module alu_74181_subset(
    input [3:0] A,  // Operand inputs
    input [3:0] B,  // Operand inputs
    input [3:0] S,  // Function selection inputs
    input M,        // Mode control input
    output reg[3:0] F   // Function outputs
    );

always @ (A, B, S, M)

// TODO

endmodule
