package tlight_package;
  typedef enum logic [2:0]{
    RED = 3'b100, 
    YELLOW = 3'b010, 
    GREEN = 3'b001} tlight_control_t;
endpackage