//
// Four-digits decimal counter
// 

module decimal_counter(
  input clock, reset,
  output logic [3:0][3:0] digits);

// TODO

endmodule